magic
tech gf180mcuD
magscale 1 10
timestamp 1765203931
<< nwell >>
rect -86 352 3222 870
<< pwell >>
rect -86 -86 3222 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 716 68 836 232
rect 940 68 1060 232
rect 1388 68 1508 232
rect 1759 68 1879 232
rect 2207 68 2327 232
rect 2575 68 2695 232
rect 2799 68 2919 232
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 716 472 816 716
rect 940 472 1040 716
rect 1164 472 1264 716
rect 1759 472 1859 716
rect 1983 472 2083 716
rect 2575 472 2675 716
rect 2799 472 2899 716
<< mvndiff >>
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 127 348 232
rect 244 81 273 127
rect 319 81 348 127
rect 244 68 348 81
rect 468 218 556 232
rect 468 172 497 218
rect 543 172 556 218
rect 468 68 556 172
rect 628 218 716 232
rect 628 172 641 218
rect 687 172 716 218
rect 628 68 716 172
rect 836 127 940 232
rect 836 81 865 127
rect 911 81 940 127
rect 836 68 940 81
rect 1060 68 1388 232
rect 1508 219 1596 232
rect 1508 173 1537 219
rect 1583 173 1596 219
rect 1508 68 1596 173
rect 1668 127 1759 232
rect 1668 81 1684 127
rect 1730 81 1759 127
rect 1668 68 1759 81
rect 1879 68 2207 232
rect 2327 218 2415 232
rect 2327 172 2356 218
rect 2402 172 2415 218
rect 2327 68 2415 172
rect 2487 127 2575 232
rect 2487 81 2500 127
rect 2546 81 2575 127
rect 2487 68 2575 81
rect 2695 219 2799 232
rect 2695 173 2724 219
rect 2770 173 2799 219
rect 2695 68 2799 173
rect 2919 127 3007 232
rect 2919 81 2948 127
rect 2994 81 3007 127
rect 2919 68 3007 81
<< mvpdiff >>
rect 36 575 124 716
rect 36 529 49 575
rect 95 529 124 575
rect 36 472 124 529
rect 224 703 348 716
rect 224 657 253 703
rect 299 657 348 703
rect 224 472 348 657
rect 448 531 556 716
rect 448 485 497 531
rect 543 485 556 531
rect 448 472 556 485
rect 628 531 716 716
rect 628 485 641 531
rect 687 485 716 531
rect 628 472 716 485
rect 816 703 940 716
rect 816 657 854 703
rect 900 657 940 703
rect 816 472 940 657
rect 1040 472 1164 716
rect 1264 531 1596 716
rect 1264 485 1537 531
rect 1583 485 1596 531
rect 1264 472 1596 485
rect 1668 703 1759 716
rect 1668 657 1681 703
rect 1727 657 1759 703
rect 1668 472 1759 657
rect 1859 472 1983 716
rect 2083 531 2415 716
rect 2083 485 2356 531
rect 2402 485 2415 531
rect 2083 472 2415 485
rect 2487 703 2575 716
rect 2487 657 2500 703
rect 2546 657 2575 703
rect 2487 472 2575 657
rect 2675 667 2799 716
rect 2675 485 2724 667
rect 2770 485 2799 667
rect 2675 472 2799 485
rect 2899 703 2987 716
rect 2899 657 2928 703
rect 2974 657 2987 703
rect 2899 472 2987 657
<< mvndiffc >>
rect 49 173 95 219
rect 273 81 319 127
rect 497 172 543 218
rect 641 172 687 218
rect 865 81 911 127
rect 1537 173 1583 219
rect 1684 81 1730 127
rect 2356 172 2402 218
rect 2500 81 2546 127
rect 2724 173 2770 219
rect 2948 81 2994 127
<< mvpdiffc >>
rect 49 529 95 575
rect 253 657 299 703
rect 497 485 543 531
rect 641 485 687 531
rect 854 657 900 703
rect 1537 485 1583 531
rect 1681 657 1727 703
rect 2356 485 2402 531
rect 2500 657 2546 703
rect 2724 485 2770 667
rect 2928 657 2974 703
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 716 716 816 760
rect 940 716 1040 760
rect 1164 716 1264 760
rect 1759 716 1859 760
rect 1983 716 2083 760
rect 2575 716 2675 760
rect 2799 716 2899 760
rect 124 439 224 472
rect 124 276 141 439
rect 187 276 224 439
rect 348 428 448 472
rect 348 382 361 428
rect 407 382 448 428
rect 348 349 448 382
rect 716 349 816 472
rect 940 349 1040 472
rect 1164 410 1264 472
rect 1164 364 1186 410
rect 1232 364 1264 410
rect 1164 349 1264 364
rect 1759 375 1859 472
rect 348 325 468 349
rect 348 279 361 325
rect 407 279 468 325
rect 124 232 244 276
rect 348 232 468 279
rect 716 346 836 349
rect 716 300 752 346
rect 798 300 836 346
rect 716 232 836 300
rect 940 311 1060 349
rect 940 265 953 311
rect 999 265 1060 311
rect 940 232 1060 265
rect 1388 333 1508 349
rect 1388 287 1423 333
rect 1469 287 1508 333
rect 1388 232 1508 287
rect 1759 329 1778 375
rect 1824 349 1859 375
rect 1983 408 2083 472
rect 1983 362 2008 408
rect 2054 362 2083 408
rect 1983 349 2083 362
rect 2575 393 2675 472
rect 2799 393 2899 472
rect 2575 385 2919 393
rect 1824 329 1879 349
rect 1759 232 1879 329
rect 2207 336 2327 349
rect 2207 290 2241 336
rect 2287 290 2327 336
rect 2207 232 2327 290
rect 2575 339 2593 385
rect 2639 339 2919 385
rect 2575 328 2919 339
rect 2575 232 2695 328
rect 2799 232 2919 328
rect 124 24 244 68
rect 348 24 468 68
rect 716 24 836 68
rect 940 24 1060 68
rect 1388 24 1508 68
rect 1759 24 1879 68
rect 2207 24 2327 68
rect 2575 24 2695 68
rect 2799 24 2919 68
<< polycontact >>
rect 141 276 187 439
rect 361 382 407 428
rect 1186 364 1232 410
rect 361 279 407 325
rect 752 300 798 346
rect 953 265 999 311
rect 1423 287 1469 333
rect 1778 329 1824 375
rect 2008 362 2054 408
rect 2241 290 2287 336
rect 2593 339 2639 385
<< metal1 >>
rect 0 724 3136 844
rect 253 703 299 724
rect 253 646 299 657
rect 854 703 900 724
rect 854 646 900 657
rect 1681 703 1727 724
rect 1681 646 1727 657
rect 2500 703 2546 724
rect 2928 703 2974 724
rect 2500 646 2546 657
rect 2722 667 2776 678
rect 493 629 551 641
rect 49 575 95 590
rect 493 577 497 629
rect 549 577 551 629
rect 95 529 407 575
rect 493 565 551 577
rect 1664 585 2271 591
rect 49 518 95 529
rect 122 439 222 466
rect 122 276 141 439
rect 187 276 222 439
rect 361 428 407 529
rect 361 325 407 382
rect 361 255 407 279
rect 497 531 543 565
rect 341 243 415 255
rect 49 230 95 232
rect 341 230 351 243
rect 49 219 351 230
rect 95 191 351 219
rect 403 191 415 243
rect 95 184 415 191
rect 497 218 543 485
rect 49 162 95 173
rect 497 161 543 172
rect 641 531 687 542
rect 641 230 687 485
rect 1537 531 1583 542
rect 1664 533 1676 585
rect 1728 545 2271 585
rect 1728 533 1740 545
rect 1664 530 1740 533
rect 733 346 834 467
rect 1164 413 1264 424
rect 1164 361 1186 413
rect 1238 361 1264 413
rect 1164 349 1264 361
rect 1537 375 1583 485
rect 1986 408 2079 424
rect 733 300 752 346
rect 798 300 834 346
rect 1398 335 1491 349
rect 733 276 834 300
rect 953 311 999 322
rect 1398 283 1420 335
rect 1472 283 1491 335
rect 1398 274 1491 283
rect 1537 329 1778 375
rect 1824 329 1840 375
rect 1986 362 2008 408
rect 2054 362 2079 408
rect 1986 349 2079 362
rect 2225 349 2271 545
rect 2356 531 2402 542
rect 2356 393 2402 485
rect 2722 485 2724 667
rect 2770 485 2776 667
rect 2928 646 2974 657
rect 2356 385 2650 393
rect 953 230 999 265
rect 641 218 999 230
rect 687 184 999 218
rect 1537 219 1583 329
rect 641 161 687 172
rect 1537 161 1583 173
rect 1776 170 1845 182
rect 273 127 319 138
rect 273 60 319 81
rect 865 127 911 138
rect 865 60 911 81
rect 1684 127 1730 138
rect 1776 118 1781 170
rect 1833 157 1845 170
rect 2005 157 2051 349
rect 2219 336 2307 349
rect 2219 290 2241 336
rect 2287 290 2307 336
rect 2219 274 2307 290
rect 2356 339 2593 385
rect 2639 339 2650 385
rect 2356 328 2650 339
rect 2356 218 2402 328
rect 2356 161 2402 172
rect 2722 219 2776 485
rect 2722 173 2724 219
rect 2770 173 2776 219
rect 2722 158 2776 173
rect 1833 118 2051 157
rect 1776 111 2051 118
rect 2500 127 2546 138
rect 1776 106 1847 111
rect 1684 60 1730 81
rect 2500 60 2546 81
rect 2948 127 2994 138
rect 2948 60 2994 81
rect 0 -60 3136 60
<< via1 >>
rect 497 577 549 629
rect 351 191 403 243
rect 1676 533 1728 585
rect 1186 410 1238 413
rect 1186 364 1232 410
rect 1232 364 1238 410
rect 1186 361 1238 364
rect 1420 333 1472 335
rect 1420 287 1423 333
rect 1423 287 1469 333
rect 1469 287 1472 333
rect 1420 283 1472 287
rect 1781 118 1833 170
<< metal2 >>
rect 493 629 551 641
rect 493 577 497 629
rect 549 622 551 629
rect 549 589 1239 622
rect 549 585 1740 589
rect 549 577 1676 585
rect 493 566 1676 577
rect 493 565 551 566
rect 1183 533 1676 566
rect 1728 533 1740 585
rect 1183 425 1239 533
rect 1672 531 1740 533
rect 1183 413 1240 425
rect 1183 361 1186 413
rect 1238 361 1240 413
rect 1183 349 1240 361
rect 1417 335 1474 347
rect 1417 283 1420 335
rect 1472 283 1474 335
rect 1417 280 1474 283
rect 347 243 406 255
rect 347 191 351 243
rect 403 191 406 243
rect 347 187 406 191
rect 348 162 406 187
rect 1417 162 1473 280
rect 1769 170 1846 172
rect 1769 162 1781 170
rect 348 118 1781 162
rect 1833 118 1846 170
rect 348 106 1846 118
<< labels >>
flabel metal1 s 0 724 3136 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 3136 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 122 276 222 466 0 FreeSans 400 0 0 0 CLK
port 7 nsew clock input
flabel metal1 733 276 834 467 0 FreeSans 200 0 0 0 D
port 5 nsew signal input
flabel metal1 2722 158 2776 678 0 FreeSans 200 0 0 0 Q
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 3136 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -40 3152 352
string MASKHINTS_PPLUS -16 352 3152 824
<< end >>
