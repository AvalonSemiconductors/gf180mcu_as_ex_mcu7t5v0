VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t5v0__trans_2
  CLASS core ;
  FOREIGN gf180mcu_as_sc_mcu7t5v0__trans_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.330 0.810 1.630 2.930 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.978400 ;
    PORT
      LAYER Metal1 ;
        RECT 0.180 0.810 0.475 3.390 ;
    END
    PORT
      LAYER Pwell ;
        RECT 2.375 0.810 2.770 1.150 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 2.375 1.150 2.670 3.390 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0.475 3.160 2.375 3.390 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 3.360 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 0.050 3.670 0.550 4.170 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.050 -0.250 0.550 0.250 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 3.360 0.300 ;
    END
  END VSS
  PIN ENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Nwell ;
        RECT 0.705 1.910 0.975 2.930 ;
    END
  END ENB
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Pwell ;
        RECT 0.710 0.530 0.985 1.610 ;
    END
  END EN
  OBS
      LAYER Nwell ;
        RECT -0.430 4.170 3.790 4.350 ;
        RECT -0.430 3.670 0.050 4.170 ;
        RECT 0.550 3.670 3.790 4.170 ;
        RECT -0.430 2.930 3.790 3.670 ;
        RECT -0.430 1.910 0.705 2.930 ;
        RECT 0.975 1.910 3.790 2.930 ;
        RECT -0.430 1.760 3.790 1.910 ;
      LAYER Pwell ;
        RECT -0.430 1.610 3.790 1.760 ;
        RECT -0.430 0.530 0.710 1.610 ;
      LAYER Nwell ;
        RECT 0.710 1.150 0.985 1.310 ;
      LAYER Pwell ;
        RECT 0.985 1.150 3.790 1.610 ;
      LAYER Nwell ;
        RECT 0.710 0.810 2.770 1.150 ;
      LAYER Pwell ;
        RECT 2.770 0.810 3.790 1.150 ;
      LAYER Nwell ;
        RECT 0.710 0.530 0.985 0.810 ;
      LAYER Pwell ;
        RECT 0.985 0.530 3.790 0.810 ;
        RECT -0.430 0.250 3.790 0.530 ;
        RECT -0.430 -0.250 0.050 0.250 ;
      LAYER Nwell ;
        RECT 0.050 0.000 0.550 0.250 ;
      LAYER Pwell ;
        RECT 0.550 -0.250 3.790 0.250 ;
        RECT -0.430 -0.430 3.790 -0.250 ;
      LAYER Metal1 ;
        RECT 0.775 0.600 1.030 2.860 ;
        RECT 1.930 0.850 2.075 2.860 ;
        RECT 1.930 0.600 2.770 0.850 ;
  END
END gf180mcu_as_sc_mcu7t5v0__trans_2
END LIBRARY

