magic
tech gf180mcuD
magscale 1 10
timestamp 1757970249
<< nwell >>
rect -86 352 3782 870
<< pwell >>
rect -86 -86 3782 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 716 68 836 232
rect 996 68 1116 232
rect 1396 68 1516 232
rect 1564 68 1684 232
rect 1788 68 1908 232
rect 2012 68 2132 232
rect 2324 68 2444 232
rect 2554 68 2674 232
rect 2778 68 2898 232
rect 3148 68 3268 232
rect 3372 68 3492 232
<< mvpmos >>
rect 124 472 224 716
rect 348 472 448 716
rect 848 472 948 716
rect 996 472 1096 716
rect 1220 472 1320 716
rect 1564 472 1664 716
rect 1788 472 1888 716
rect 2120 472 2220 716
rect 2406 472 2506 716
rect 2554 472 2654 716
rect 2778 472 2878 716
rect 3148 472 3248 716
rect 3372 472 3472 716
<< mvndiff >>
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 127 348 232
rect 244 81 273 127
rect 319 81 348 127
rect 244 68 348 81
rect 468 218 556 232
rect 468 172 497 218
rect 543 172 556 218
rect 468 68 556 172
rect 628 127 716 232
rect 628 81 641 127
rect 687 81 716 127
rect 628 68 716 81
rect 836 68 996 232
rect 1116 219 1396 232
rect 1116 173 1145 219
rect 1191 173 1396 219
rect 1116 68 1396 173
rect 1516 68 1564 232
rect 1684 127 1788 232
rect 1684 81 1713 127
rect 1759 81 1788 127
rect 1684 68 1788 81
rect 1908 219 2012 232
rect 1908 173 1937 219
rect 1983 173 2012 219
rect 1908 68 2012 173
rect 2132 219 2324 232
rect 2132 173 2249 219
rect 2295 173 2324 219
rect 2132 68 2324 173
rect 2444 68 2554 232
rect 2674 127 2778 232
rect 2674 81 2703 127
rect 2749 81 2778 127
rect 2674 68 2778 81
rect 2898 219 2986 232
rect 2898 173 2927 219
rect 2973 173 2986 219
rect 2898 68 2986 173
rect 3058 127 3148 232
rect 3058 81 3073 127
rect 3119 81 3148 127
rect 3058 68 3148 81
rect 3268 219 3372 232
rect 3268 173 3297 219
rect 3343 173 3372 219
rect 3268 68 3372 173
rect 3492 127 3580 232
rect 3492 81 3521 127
rect 3567 81 3580 127
rect 3492 68 3580 81
<< mvpdiff >>
rect 36 575 124 716
rect 36 529 49 575
rect 95 529 124 575
rect 36 472 124 529
rect 224 703 348 716
rect 224 657 253 703
rect 299 657 348 703
rect 224 472 348 657
rect 448 531 556 716
rect 448 485 497 531
rect 543 485 556 531
rect 448 472 556 485
rect 628 703 848 716
rect 628 656 760 703
rect 806 656 848 703
rect 628 472 848 656
rect 948 472 996 716
rect 1096 531 1220 716
rect 1096 485 1145 531
rect 1191 485 1220 531
rect 1096 472 1220 485
rect 1320 472 1564 716
rect 1664 702 1788 716
rect 1664 656 1693 702
rect 1739 656 1788 702
rect 1664 472 1788 656
rect 1888 531 2120 716
rect 1888 485 1937 531
rect 1983 485 2120 531
rect 1888 472 2120 485
rect 2220 531 2406 716
rect 2220 485 2249 531
rect 2295 485 2406 531
rect 2220 472 2406 485
rect 2506 472 2554 716
rect 2654 703 2778 716
rect 2654 657 2683 703
rect 2729 657 2778 703
rect 2654 472 2778 657
rect 2878 667 2986 716
rect 2878 485 2927 667
rect 2973 485 2986 667
rect 2878 472 2986 485
rect 3058 703 3148 716
rect 3058 485 3071 703
rect 3117 485 3148 703
rect 3058 472 3148 485
rect 3248 667 3372 716
rect 3248 485 3297 667
rect 3343 485 3372 667
rect 3248 472 3372 485
rect 3472 703 3562 716
rect 3472 485 3503 703
rect 3549 485 3562 703
rect 3472 472 3562 485
<< mvndiffc >>
rect 49 173 95 219
rect 273 81 319 127
rect 497 172 543 218
rect 641 81 687 127
rect 1145 173 1191 219
rect 1713 81 1759 127
rect 1937 173 1983 219
rect 2249 173 2295 219
rect 2703 81 2749 127
rect 2927 173 2973 219
rect 3073 81 3119 127
rect 3297 173 3343 219
rect 3521 81 3567 127
<< mvpdiffc >>
rect 49 529 95 575
rect 253 657 299 703
rect 497 485 543 531
rect 760 656 806 703
rect 1145 485 1191 531
rect 1693 656 1739 702
rect 1937 485 1983 531
rect 2249 485 2295 531
rect 2683 657 2729 703
rect 2927 485 2973 667
rect 3071 485 3117 703
rect 3297 485 3343 667
rect 3503 485 3549 703
<< polysilicon >>
rect 124 716 224 760
rect 348 716 448 760
rect 848 716 948 760
rect 996 716 1096 760
rect 1220 716 1320 760
rect 1564 716 1664 760
rect 1788 716 1888 760
rect 2120 716 2220 760
rect 2406 716 2506 760
rect 2554 716 2654 760
rect 2778 716 2878 760
rect 3148 716 3248 760
rect 3372 716 3472 760
rect 124 439 224 472
rect 124 276 141 439
rect 187 276 224 439
rect 348 428 448 472
rect 348 382 361 428
rect 407 382 448 428
rect 848 439 948 472
rect 848 397 889 439
rect 348 349 448 382
rect 876 393 889 397
rect 935 393 948 439
rect 876 364 948 393
rect 996 434 1096 472
rect 996 388 1009 434
rect 1056 388 1096 434
rect 1220 439 1320 472
rect 1220 428 1250 439
rect 348 325 829 349
rect 348 279 361 325
rect 407 311 829 325
rect 996 331 1096 388
rect 1237 392 1250 428
rect 1298 392 1320 439
rect 1237 379 1320 392
rect 407 292 836 311
rect 407 279 468 292
rect 124 232 244 276
rect 348 232 468 279
rect 716 232 836 292
rect 996 285 1009 331
rect 1056 285 1096 331
rect 996 276 1096 285
rect 1433 336 1516 356
rect 1433 289 1451 336
rect 1499 289 1516 336
rect 1433 276 1516 289
rect 996 232 1116 276
rect 1396 232 1516 276
rect 1564 354 1664 472
rect 1788 412 1888 472
rect 2120 439 2220 472
rect 2120 428 2152 439
rect 1564 307 1577 354
rect 1625 307 1664 354
rect 1774 399 1888 412
rect 1774 352 1790 399
rect 1838 352 1888 399
rect 2139 393 2152 428
rect 2198 393 2220 439
rect 2406 439 2506 472
rect 2406 428 2447 439
rect 2139 380 2220 393
rect 2434 393 2447 428
rect 2493 393 2506 439
rect 2434 380 2506 393
rect 2554 390 2654 472
rect 1774 339 1888 352
rect 2155 367 2220 380
rect 1564 289 1664 307
rect 1564 232 1684 289
rect 1788 276 1888 339
rect 2029 327 2101 348
rect 2029 281 2042 327
rect 2088 281 2101 327
rect 2155 319 2376 367
rect 2029 276 2101 281
rect 2324 276 2376 319
rect 2554 344 2595 390
rect 2641 344 2654 390
rect 2554 276 2654 344
rect 2778 317 2878 472
rect 3148 390 3248 472
rect 3372 390 3472 472
rect 1788 232 1908 276
rect 2012 232 2132 276
rect 2324 232 2444 276
rect 2554 232 2674 276
rect 2778 271 2792 317
rect 2838 277 2878 317
rect 2982 374 3472 390
rect 2982 328 2995 374
rect 3041 328 3472 374
rect 2982 313 3472 328
rect 2838 271 2898 277
rect 2778 232 2898 271
rect 3148 232 3268 313
rect 3372 280 3472 313
rect 3372 232 3492 280
rect 124 24 244 68
rect 348 24 468 68
rect 716 24 836 68
rect 996 24 1116 68
rect 1396 24 1516 68
rect 1564 24 1684 68
rect 1788 24 1908 68
rect 2012 24 2132 68
rect 2324 24 2444 68
rect 2554 24 2674 68
rect 2778 24 2898 68
rect 3148 24 3268 68
rect 3372 24 3492 68
<< polycontact >>
rect 141 276 187 439
rect 361 382 407 428
rect 889 393 935 439
rect 1009 388 1056 434
rect 361 279 407 325
rect 1250 392 1298 439
rect 1009 285 1056 331
rect 1451 289 1499 336
rect 1577 307 1625 354
rect 1790 352 1838 399
rect 2152 393 2198 439
rect 2447 393 2493 439
rect 2042 281 2088 327
rect 2595 344 2641 390
rect 2792 271 2838 317
rect 2995 328 3041 374
<< metal1 >>
rect 0 724 3696 844
rect 253 703 299 724
rect 253 646 299 657
rect 760 703 806 724
rect 760 645 806 656
rect 1693 702 1739 724
rect 1693 645 1739 656
rect 2683 703 2729 724
rect 3071 703 3117 724
rect 2683 646 2729 657
rect 2927 667 2973 678
rect 49 575 95 590
rect 353 588 665 634
rect 353 575 407 588
rect 95 529 407 575
rect 617 581 665 588
rect 1053 598 1644 634
rect 1799 604 1875 605
rect 1799 598 1811 604
rect 1053 588 1811 598
rect 1053 581 1099 588
rect 49 518 95 529
rect 122 439 222 466
rect 122 276 141 439
rect 187 276 222 439
rect 361 428 407 529
rect 361 325 407 382
rect 49 230 95 232
rect 361 230 407 279
rect 49 219 407 230
rect 95 184 407 219
rect 497 531 543 542
rect 617 535 1099 581
rect 497 449 543 485
rect 1145 531 1191 542
rect 876 449 935 450
rect 497 439 935 449
rect 497 393 889 439
rect 497 390 935 393
rect 497 218 543 390
rect 876 382 935 390
rect 49 162 95 173
rect 497 161 543 172
rect 887 152 935 382
rect 996 434 1096 463
rect 996 388 1009 434
rect 1056 388 1096 434
rect 996 331 1096 388
rect 996 285 1009 331
rect 1056 285 1096 331
rect 996 273 1096 285
rect 1145 346 1191 485
rect 1237 445 1298 588
rect 1593 552 1811 588
rect 1863 552 1875 604
rect 2044 588 2499 634
rect 1937 531 1983 542
rect 1237 439 1309 445
rect 1237 392 1250 439
rect 1298 392 1309 439
rect 1355 413 1839 460
rect 1355 346 1403 413
rect 1790 399 1839 413
rect 1145 300 1403 346
rect 1449 340 1522 356
rect 1145 219 1191 300
rect 1449 288 1451 340
rect 1503 288 1522 340
rect 1449 276 1522 288
rect 1568 354 1632 362
rect 1568 307 1577 354
rect 1625 307 1632 354
rect 1838 352 1839 399
rect 1790 341 1839 352
rect 1568 231 1632 307
rect 1937 231 1983 485
rect 2044 352 2090 588
rect 2249 531 2295 542
rect 2139 447 2203 459
rect 2139 395 2143 447
rect 2195 439 2203 447
rect 2139 393 2152 395
rect 2198 393 2203 439
rect 2139 368 2203 393
rect 2029 340 2090 352
rect 2029 288 2031 340
rect 2083 327 2090 340
rect 2029 281 2042 288
rect 2088 281 2090 327
rect 2029 251 2090 281
rect 1568 219 1983 231
rect 1568 185 1937 219
rect 1145 162 1191 173
rect 1937 162 1983 173
rect 2249 236 2295 485
rect 2436 439 2499 588
rect 2927 467 2973 485
rect 2436 393 2447 439
rect 2493 393 2499 439
rect 2436 382 2499 393
rect 2595 421 2973 467
rect 3503 703 3549 724
rect 3071 452 3117 485
rect 3284 667 3361 678
rect 3284 485 3297 667
rect 3343 485 3361 667
rect 2595 390 2641 421
rect 2595 332 2641 344
rect 2927 374 2973 421
rect 2927 328 2995 374
rect 3041 328 3052 374
rect 2791 317 2840 328
rect 2791 271 2792 317
rect 2838 271 2840 317
rect 2791 236 2840 271
rect 2249 219 2840 236
rect 2295 184 2840 219
rect 2927 219 2973 328
rect 2249 162 2295 173
rect 2927 162 2973 173
rect 3284 219 3361 485
rect 3503 458 3549 485
rect 3284 173 3297 219
rect 3343 173 3361 219
rect 1006 152 1018 160
rect 273 127 319 138
rect 273 60 319 81
rect 641 127 687 138
rect 887 108 1018 152
rect 1070 108 1082 160
rect 3284 147 3361 173
rect 887 106 1082 108
rect 1713 127 1759 138
rect 641 60 687 81
rect 1713 60 1759 81
rect 2703 127 2749 138
rect 2703 60 2749 81
rect 3073 127 3119 138
rect 3073 60 3119 81
rect 3521 127 3567 138
rect 3521 60 3567 81
rect 0 -60 3696 60
<< via1 >>
rect 1811 552 1863 604
rect 1451 336 1503 340
rect 1451 289 1499 336
rect 1499 289 1503 336
rect 1451 288 1503 289
rect 2143 439 2195 447
rect 2143 395 2152 439
rect 2152 395 2195 439
rect 2031 327 2083 340
rect 2031 288 2042 327
rect 2042 288 2083 327
rect 1018 108 1070 160
<< metal2 >>
rect 1799 605 1875 607
rect 1799 604 2199 605
rect 1799 552 1811 604
rect 1863 552 2199 604
rect 1799 549 2199 552
rect 2139 447 2199 549
rect 2139 395 2143 447
rect 2195 395 2199 447
rect 2139 383 2199 395
rect 1449 342 1505 352
rect 1449 340 2095 342
rect 1449 288 1451 340
rect 1503 288 2031 340
rect 2083 288 2095 340
rect 1449 286 2095 288
rect 1449 162 1505 286
rect 1006 160 1505 162
rect 1006 108 1018 160
rect 1070 108 1505 160
rect 1006 106 1505 108
<< labels >>
flabel metal1 s 0 724 3696 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 3696 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 3284 147 3361 678 0 FreeSans 400 0 0 0 Q
port 5 nsew signal output
flabel metal1 996 273 1096 463 0 FreeSans 400 0 0 0 D
port 6 nsew signal input
flabel metal1 122 276 222 466 0 FreeSans 400 0 0 0 CLK
port 7 nsew clock input
<< properties >>
string FIXED_BBOX 0 0 3696 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string MASKHINTS_NPLUS -16 -46 3712 352
string MASKHINTS_PPLUS -16 352 3712 830
<< end >>
