VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_as_sc_mcu7t5v0__trans_1
  CLASS core ;
  FOREIGN gf180mcu_as_sc_mcu7t5v0__trans_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.240 BY 3.920 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.080800 ;
    PORT
      LAYER Metal1 ;
        RECT 1.330 0.810 1.630 3.390 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal1 ;
        RECT 0.180 0.810 0.475 3.390 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 3.620 2.240 4.220 ;
    END
  END VDD
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Nwell ;
        RECT 0.050 3.670 0.550 4.170 ;
    END
  END VNW
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Pwell ;
        RECT 0.050 -0.250 0.550 0.250 ;
    END
  END VPW
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.300 2.240 0.300 ;
    END
  END VSS
  PIN ENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.610000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.705 1.910 0.975 3.235 ;
    END
  END ENB
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.710 0.530 0.985 1.610 ;
    END
  END EN
  OBS
      LAYER Nwell ;
        RECT -0.430 4.170 2.670 4.350 ;
        RECT -0.430 3.670 0.050 4.170 ;
        RECT 0.550 3.670 2.670 4.170 ;
        RECT -0.430 1.760 2.670 3.670 ;
      LAYER Pwell ;
        RECT -0.430 0.250 2.670 1.760 ;
        RECT -0.430 -0.250 0.050 0.250 ;
      LAYER Nwell ;
        RECT 0.050 0.000 0.550 0.250 ;
      LAYER Pwell ;
        RECT 0.550 -0.250 2.670 0.250 ;
        RECT -0.430 -0.430 2.670 -0.250 ;
  END
END gf180mcu_as_sc_mcu7t5v0__trans_1
END LIBRARY

