magic
tech gf180mcuD
magscale 1 10
timestamp 1756916228
<< nwell >>
rect -86 377 6806 870
rect -86 352 1085 377
rect 1336 352 4109 377
rect 4360 352 6806 377
<< pwell >>
rect 1085 352 1336 377
rect 4109 352 4360 377
rect -86 -86 6806 352
<< mvnmos >>
rect 116 68 236 232
rect 341 68 461 232
rect 828 159 948 231
rect 996 159 1116 231
rect 1320 159 1440 231
rect 1488 159 1608 231
rect 1800 159 1920 231
rect 2024 159 2144 231
rect 2248 159 2368 231
rect 2416 159 2536 231
rect 2684 151 2804 231
rect 3072 68 3192 232
rect 3296 68 3416 232
rect 3852 159 3972 231
rect 4020 159 4140 231
rect 4344 159 4464 231
rect 4512 159 4632 231
rect 4824 159 4944 231
rect 5048 159 5168 231
rect 5272 159 5392 231
rect 5440 159 5560 231
rect 5708 151 5828 231
rect 6096 68 6216 232
rect 6320 68 6440 232
<< mvpmos >>
rect 122 508 222 716
rect 346 508 446 716
rect 892 527 992 599
rect 1052 527 1152 599
rect 1360 527 1460 599
rect 1508 527 1608 599
rect 1724 527 1824 599
rect 2023 527 2123 599
rect 2308 527 2408 599
rect 2464 527 2564 599
rect 2712 527 2812 687
rect 3060 472 3160 716
rect 3264 472 3364 716
rect 3916 527 4016 599
rect 4076 527 4176 599
rect 4384 527 4484 599
rect 4532 527 4632 599
rect 4748 527 4848 599
rect 5047 527 5147 599
rect 5332 527 5432 599
rect 5488 527 5588 599
rect 5736 527 5836 687
rect 6084 472 6184 716
rect 6288 472 6388 716
<< mvndiff >>
rect 28 192 116 232
rect 28 146 41 192
rect 87 146 116 192
rect 28 68 116 146
rect 236 143 341 232
rect 236 97 266 143
rect 312 97 341 143
rect 236 68 341 97
rect 461 219 623 232
rect 1176 244 1248 257
rect 1176 231 1189 244
rect 461 173 490 219
rect 536 173 623 219
rect 461 68 623 173
rect 696 159 828 231
rect 948 159 996 231
rect 1116 198 1189 231
rect 1235 231 1248 244
rect 1235 198 1320 231
rect 1116 159 1320 198
rect 1440 159 1488 231
rect 1608 159 1800 231
rect 1920 218 2024 231
rect 1920 172 1949 218
rect 1995 172 2024 218
rect 1920 159 2024 172
rect 2144 218 2248 231
rect 2144 172 2173 218
rect 2219 172 2248 218
rect 2144 159 2248 172
rect 2368 159 2416 231
rect 2536 210 2684 231
rect 2536 164 2609 210
rect 2655 164 2684 210
rect 2536 159 2684 164
rect 696 143 768 159
rect 696 97 709 143
rect 755 97 768 143
rect 1668 117 1740 159
rect 696 79 768 97
rect 1668 71 1681 117
rect 1727 71 1740 117
rect 2596 151 2684 159
rect 2804 210 2892 231
rect 2804 164 2833 210
rect 2879 164 2892 210
rect 2804 151 2892 164
rect 2984 167 3072 232
rect 1668 58 1740 71
rect 2984 121 2997 167
rect 3043 121 3072 167
rect 2984 68 3072 121
rect 3192 167 3296 232
rect 3192 121 3221 167
rect 3267 121 3296 167
rect 3192 68 3296 121
rect 3416 158 3616 232
rect 4200 244 4272 257
rect 4200 231 4213 244
rect 3416 112 3445 158
rect 3491 112 3616 158
rect 3416 68 3616 112
rect 3720 159 3852 231
rect 3972 159 4020 231
rect 4140 198 4213 231
rect 4259 231 4272 244
rect 4259 198 4344 231
rect 4140 159 4344 198
rect 4464 159 4512 231
rect 4632 159 4824 231
rect 4944 218 5048 231
rect 4944 172 4973 218
rect 5019 172 5048 218
rect 4944 159 5048 172
rect 5168 218 5272 231
rect 5168 172 5197 218
rect 5243 172 5272 218
rect 5168 159 5272 172
rect 5392 159 5440 231
rect 5560 210 5708 231
rect 5560 164 5633 210
rect 5679 164 5708 210
rect 5560 159 5708 164
rect 3720 143 3792 159
rect 3720 97 3733 143
rect 3779 97 3792 143
rect 4692 117 4764 159
rect 3720 79 3792 97
rect 4692 71 4705 117
rect 4751 71 4764 117
rect 5620 151 5708 159
rect 5828 210 5916 231
rect 5828 164 5857 210
rect 5903 164 5916 210
rect 5828 151 5916 164
rect 6008 167 6096 232
rect 4692 58 4764 71
rect 6008 121 6021 167
rect 6067 121 6096 167
rect 6008 68 6096 121
rect 6216 167 6320 232
rect 6216 121 6245 167
rect 6291 121 6320 167
rect 6216 68 6320 121
rect 6440 158 6640 232
rect 6440 112 6469 158
rect 6515 112 6640 158
rect 6440 68 6640 112
<< mvpdiff >>
rect 34 622 122 716
rect 34 576 47 622
rect 93 576 122 622
rect 34 508 122 576
rect 222 697 346 716
rect 222 651 251 697
rect 297 651 346 697
rect 222 508 346 651
rect 446 586 638 716
rect 446 540 490 586
rect 536 540 638 586
rect 446 508 638 540
rect 760 694 832 720
rect 760 648 773 694
rect 819 648 832 694
rect 760 599 832 648
rect 2972 689 3060 716
rect 2624 599 2712 687
rect 760 527 892 599
rect 992 527 1052 599
rect 1152 586 1360 599
rect 1152 540 1245 586
rect 1291 540 1360 586
rect 1152 527 1360 540
rect 1460 527 1508 599
rect 1608 586 1724 599
rect 1608 540 1649 586
rect 1695 540 1724 586
rect 1608 527 1724 540
rect 1824 586 2023 599
rect 1824 540 1948 586
rect 1994 540 2023 586
rect 1824 527 2023 540
rect 2123 586 2308 599
rect 2123 540 2173 586
rect 2219 540 2308 586
rect 2123 527 2308 540
rect 2408 527 2464 599
rect 2564 595 2712 599
rect 2564 549 2637 595
rect 2683 549 2712 595
rect 2564 527 2712 549
rect 2812 595 2900 687
rect 2812 549 2841 595
rect 2887 549 2900 595
rect 2812 527 2900 549
rect 2972 549 2985 689
rect 3031 549 3060 689
rect 2972 472 3060 549
rect 3160 595 3264 716
rect 3160 549 3189 595
rect 3235 549 3264 595
rect 3160 472 3264 549
rect 3364 685 3584 716
rect 3364 545 3402 685
rect 3448 545 3584 685
rect 3364 472 3584 545
rect 3784 694 3856 720
rect 3784 648 3797 694
rect 3843 648 3856 694
rect 3784 599 3856 648
rect 5996 689 6084 716
rect 5648 599 5736 687
rect 3784 527 3916 599
rect 4016 527 4076 599
rect 4176 586 4384 599
rect 4176 540 4269 586
rect 4315 540 4384 586
rect 4176 527 4384 540
rect 4484 527 4532 599
rect 4632 586 4748 599
rect 4632 540 4673 586
rect 4719 540 4748 586
rect 4632 527 4748 540
rect 4848 586 5047 599
rect 4848 540 4972 586
rect 5018 540 5047 586
rect 4848 527 5047 540
rect 5147 586 5332 599
rect 5147 540 5197 586
rect 5243 540 5332 586
rect 5147 527 5332 540
rect 5432 527 5488 599
rect 5588 595 5736 599
rect 5588 549 5661 595
rect 5707 549 5736 595
rect 5588 527 5736 549
rect 5836 595 5924 687
rect 5836 549 5865 595
rect 5911 549 5924 595
rect 5836 527 5924 549
rect 5996 549 6009 689
rect 6055 549 6084 689
rect 5996 472 6084 549
rect 6184 595 6288 716
rect 6184 549 6213 595
rect 6259 549 6288 595
rect 6184 472 6288 549
rect 6388 685 6608 716
rect 6388 545 6426 685
rect 6472 545 6608 685
rect 6388 472 6608 545
<< mvndiffc >>
rect 41 146 87 192
rect 266 97 312 143
rect 490 173 536 219
rect 1189 198 1235 244
rect 1949 172 1995 218
rect 2173 172 2219 218
rect 2609 164 2655 210
rect 709 97 755 143
rect 1681 71 1727 117
rect 2833 164 2879 210
rect 2997 121 3043 167
rect 3221 121 3267 167
rect 3445 112 3491 158
rect 4213 198 4259 244
rect 4973 172 5019 218
rect 5197 172 5243 218
rect 5633 164 5679 210
rect 3733 97 3779 143
rect 4705 71 4751 117
rect 5857 164 5903 210
rect 6021 121 6067 167
rect 6245 121 6291 167
rect 6469 112 6515 158
<< mvpdiffc >>
rect 47 576 93 622
rect 251 651 297 697
rect 490 540 536 586
rect 773 648 819 694
rect 1245 540 1291 586
rect 1649 540 1695 586
rect 1948 540 1994 586
rect 2173 540 2219 586
rect 2637 549 2683 595
rect 2841 549 2887 595
rect 2985 549 3031 689
rect 3189 549 3235 595
rect 3402 545 3448 685
rect 3797 648 3843 694
rect 4269 540 4315 586
rect 4673 540 4719 586
rect 4972 540 5018 586
rect 5197 540 5243 586
rect 5661 549 5707 595
rect 5865 549 5911 595
rect 6009 549 6055 689
rect 6213 549 6259 595
rect 6426 545 6472 685
<< polysilicon >>
rect 122 716 222 760
rect 346 716 446 760
rect 1360 720 2123 760
rect 1360 678 1460 720
rect 892 599 992 672
rect 1052 599 1152 672
rect 1360 632 1373 678
rect 1419 632 1460 678
rect 1360 599 1460 632
rect 1508 599 1608 672
rect 1724 599 1824 672
rect 2023 599 2123 720
rect 2308 678 2408 691
rect 2712 687 2812 760
rect 3060 716 3160 760
rect 3264 716 3364 760
rect 4384 720 5147 760
rect 2308 632 2321 678
rect 2367 632 2408 678
rect 2308 599 2408 632
rect 2464 599 2564 643
rect 122 475 222 508
rect 122 306 149 475
rect 116 281 149 306
rect 195 306 222 475
rect 346 475 446 508
rect 346 306 371 475
rect 195 281 236 306
rect 116 232 236 281
rect 341 265 371 306
rect 417 373 446 475
rect 892 467 992 527
rect 889 455 992 467
rect 889 409 914 455
rect 960 409 992 455
rect 889 395 992 409
rect 417 364 776 373
rect 417 351 848 364
rect 417 305 789 351
rect 835 332 848 351
rect 835 305 948 332
rect 1052 324 1152 527
rect 1360 471 1460 527
rect 417 292 948 305
rect 417 265 461 292
rect 341 232 461 265
rect 828 231 948 292
rect 996 317 1152 324
rect 996 311 1116 317
rect 996 265 1038 311
rect 1084 265 1116 311
rect 996 231 1116 265
rect 1320 311 1440 324
rect 1320 265 1345 311
rect 1391 265 1440 311
rect 1508 310 1608 527
rect 1724 494 1824 527
rect 1724 448 1737 494
rect 1783 448 1824 494
rect 1724 396 1824 448
rect 2023 412 2123 527
rect 2308 483 2408 527
rect 2464 416 2564 527
rect 2712 425 2812 527
rect 4384 678 4484 720
rect 3916 599 4016 672
rect 4076 599 4176 672
rect 4384 632 4397 678
rect 4443 632 4484 678
rect 4384 599 4484 632
rect 4532 599 4632 672
rect 4748 599 4848 672
rect 5047 599 5147 720
rect 5332 678 5432 691
rect 5736 687 5836 760
rect 6084 716 6184 760
rect 6288 716 6388 760
rect 5332 632 5345 678
rect 5391 632 5432 678
rect 5332 599 5432 632
rect 5488 599 5588 643
rect 1724 356 1920 396
rect 2023 372 2288 412
rect 1508 275 1549 310
rect 1320 231 1440 265
rect 1488 264 1549 275
rect 1595 264 1608 310
rect 1488 231 1608 264
rect 1800 231 1920 356
rect 2024 310 2144 323
rect 2024 264 2056 310
rect 2102 264 2144 310
rect 2024 231 2144 264
rect 2248 275 2288 372
rect 2464 326 2536 416
rect 2464 280 2477 326
rect 2523 280 2536 326
rect 2712 379 2725 425
rect 2771 379 2812 425
rect 3060 416 3160 472
rect 2712 311 2812 379
rect 3072 394 3160 416
rect 3264 394 3364 472
rect 3916 467 4016 527
rect 3913 455 4016 467
rect 3913 409 3938 455
rect 3984 409 4016 455
rect 3913 395 4016 409
rect 3072 370 3364 394
rect 3072 357 3416 370
rect 3072 311 3085 357
rect 3131 313 3416 357
rect 3131 311 3192 313
rect 2712 288 2804 311
rect 2464 275 2536 280
rect 2248 231 2368 275
rect 2416 231 2536 275
rect 2684 231 2804 288
rect 3072 232 3192 311
rect 3296 232 3416 313
rect 3800 351 3872 364
rect 3800 305 3813 351
rect 3859 332 3872 351
rect 3859 305 3972 332
rect 4076 324 4176 527
rect 4384 471 4484 527
rect 3800 292 3972 305
rect 828 115 948 159
rect 996 115 1116 159
rect 1320 115 1440 159
rect 1488 115 1608 159
rect 1800 115 1920 159
rect 2024 115 2144 159
rect 2248 115 2368 159
rect 2416 115 2536 159
rect 116 24 236 68
rect 341 24 461 68
rect 2684 24 2804 151
rect 3852 231 3972 292
rect 4020 317 4176 324
rect 4020 311 4140 317
rect 4020 265 4062 311
rect 4108 265 4140 311
rect 4020 231 4140 265
rect 4344 311 4464 324
rect 4344 265 4369 311
rect 4415 265 4464 311
rect 4532 310 4632 527
rect 4748 494 4848 527
rect 4748 448 4761 494
rect 4807 448 4848 494
rect 4748 396 4848 448
rect 5047 412 5147 527
rect 5332 483 5432 527
rect 5488 416 5588 527
rect 5736 425 5836 527
rect 4748 356 4944 396
rect 5047 372 5312 412
rect 4532 275 4573 310
rect 4344 231 4464 265
rect 4512 264 4573 275
rect 4619 264 4632 310
rect 4512 231 4632 264
rect 4824 231 4944 356
rect 5048 310 5168 323
rect 5048 264 5080 310
rect 5126 264 5168 310
rect 5048 231 5168 264
rect 5272 275 5312 372
rect 5488 326 5560 416
rect 5488 280 5501 326
rect 5547 280 5560 326
rect 5736 379 5749 425
rect 5795 379 5836 425
rect 6084 416 6184 472
rect 5736 311 5836 379
rect 6096 394 6184 416
rect 6288 394 6388 472
rect 6096 370 6388 394
rect 6096 357 6440 370
rect 6096 311 6109 357
rect 6155 313 6440 357
rect 6155 311 6216 313
rect 5736 288 5828 311
rect 5488 275 5560 280
rect 5272 231 5392 275
rect 5440 231 5560 275
rect 5708 231 5828 288
rect 6096 232 6216 311
rect 6320 232 6440 313
rect 3852 115 3972 159
rect 4020 115 4140 159
rect 4344 115 4464 159
rect 4512 115 4632 159
rect 4824 115 4944 159
rect 5048 115 5168 159
rect 5272 115 5392 159
rect 5440 115 5560 159
rect 3072 24 3192 68
rect 3296 24 3416 68
rect 5708 24 5828 151
rect 6096 24 6216 68
rect 6320 24 6440 68
<< polycontact >>
rect 1373 632 1419 678
rect 2321 632 2367 678
rect 149 281 195 475
rect 371 265 417 475
rect 914 409 960 455
rect 789 305 835 351
rect 1038 265 1084 311
rect 1345 265 1391 311
rect 1737 448 1783 494
rect 4397 632 4443 678
rect 5345 632 5391 678
rect 1549 264 1595 310
rect 2056 264 2102 310
rect 2477 280 2523 326
rect 2725 379 2771 425
rect 3938 409 3984 455
rect 3085 311 3131 357
rect 3813 305 3859 351
rect 4062 265 4108 311
rect 4369 265 4415 311
rect 4761 448 4807 494
rect 4573 264 4619 310
rect 5080 264 5126 310
rect 5501 280 5547 326
rect 5749 379 5795 425
rect 6109 311 6155 357
<< metal1 >>
rect 0 724 6720 844
rect 251 697 297 724
rect 47 622 93 678
rect 251 637 297 651
rect 773 694 819 724
rect 773 637 819 648
rect 934 632 1368 678
rect 1420 632 1432 678
rect 93 576 417 591
rect 47 545 417 576
rect 112 475 240 499
rect 112 281 149 475
rect 195 281 240 475
rect 371 475 417 545
rect 371 235 417 265
rect 41 192 417 235
rect 87 189 417 192
rect 490 586 536 603
rect 934 558 980 632
rect 1368 614 1420 626
rect 1638 586 1706 724
rect 490 237 536 540
rect 789 512 980 558
rect 789 351 835 512
rect 789 288 835 305
rect 881 455 927 465
rect 881 409 914 455
rect 960 409 973 455
rect 881 237 927 409
rect 1026 311 1107 542
rect 1234 540 1245 586
rect 1291 540 1302 586
rect 1638 540 1649 586
rect 1695 540 1706 586
rect 1840 632 2321 678
rect 2367 632 2378 678
rect 1234 494 1302 540
rect 1026 265 1038 311
rect 1084 265 1107 311
rect 1026 242 1107 265
rect 1177 448 1737 494
rect 1783 448 1794 494
rect 1177 244 1246 448
rect 1840 402 1886 632
rect 490 219 927 237
rect 536 191 927 219
rect 1177 198 1189 244
rect 1235 198 1246 244
rect 1345 356 1886 402
rect 1937 540 1948 586
rect 1994 540 2006 586
rect 1345 311 1391 356
rect 1937 310 2006 540
rect 490 162 536 173
rect 41 135 87 146
rect 881 152 927 191
rect 1345 170 1391 265
rect 1538 264 1549 310
rect 1595 264 2006 310
rect 1938 218 2006 264
rect 2056 310 2102 632
rect 2637 595 2683 724
rect 2985 689 3031 724
rect 2056 245 2102 264
rect 2162 540 2173 586
rect 2219 540 2230 586
rect 2162 426 2230 540
rect 2637 527 2683 549
rect 2841 595 2887 606
rect 2162 425 2782 426
rect 2162 379 2725 425
rect 2771 379 2782 425
rect 1938 172 1949 218
rect 1995 172 2006 218
rect 2162 218 2230 379
rect 2841 368 2887 549
rect 3402 685 3448 724
rect 2985 527 3031 549
rect 3079 549 3189 595
rect 3235 549 3282 595
rect 3079 466 3282 549
rect 3797 694 3843 724
rect 3797 637 3843 648
rect 3946 626 3958 678
rect 4010 632 4397 678
rect 4443 632 4454 678
rect 4010 626 4022 632
rect 3946 614 4022 626
rect 3958 558 4004 614
rect 4662 586 4730 724
rect 3402 527 3448 545
rect 2841 357 3131 368
rect 2841 326 3085 357
rect 2466 280 2477 326
rect 2523 311 3085 326
rect 2523 300 3131 311
rect 2523 280 2886 300
rect 2162 172 2173 218
rect 2219 172 2230 218
rect 2609 210 2655 221
rect 1327 158 1403 170
rect 1327 152 1339 158
rect 252 97 266 143
rect 312 97 326 143
rect 252 60 326 97
rect 698 97 709 143
rect 755 97 772 143
rect 881 106 1339 152
rect 1391 106 1403 158
rect 698 60 772 97
rect 1670 71 1681 117
rect 1727 71 1738 117
rect 1670 60 1738 71
rect 2609 60 2655 164
rect 2833 210 2886 280
rect 2879 164 2886 210
rect 2833 151 2886 164
rect 2997 167 3043 178
rect 2997 60 3043 121
rect 3206 167 3282 466
rect 3813 512 4004 558
rect 3813 351 3859 512
rect 3813 288 3859 305
rect 3905 455 3951 465
rect 3905 409 3938 455
rect 3984 409 3997 455
rect 3206 121 3221 167
rect 3267 121 3282 167
rect 3206 110 3282 121
rect 3445 158 3491 178
rect 3905 162 3951 409
rect 4050 311 4131 542
rect 4258 540 4269 586
rect 4315 540 4326 586
rect 4662 540 4673 586
rect 4719 540 4730 586
rect 4864 632 5345 678
rect 5391 632 5402 678
rect 4258 494 4326 540
rect 4050 254 4062 311
rect 4108 306 4131 311
rect 4114 254 4131 306
rect 4050 242 4131 254
rect 4201 448 4761 494
rect 4807 448 4818 494
rect 4201 244 4270 448
rect 4864 402 4910 632
rect 4201 198 4213 244
rect 4259 198 4270 244
rect 4369 356 4910 402
rect 4961 540 4972 586
rect 5018 540 5030 586
rect 4369 311 4415 356
rect 4961 310 5030 540
rect 3893 158 3969 162
rect 3445 60 3491 112
rect 3722 97 3733 143
rect 3779 97 3796 143
rect 3893 106 3905 158
rect 3957 152 3969 158
rect 4369 152 4415 265
rect 4562 264 4573 310
rect 4619 264 5030 310
rect 4962 218 5030 264
rect 5080 310 5126 632
rect 5661 595 5707 724
rect 6009 689 6055 724
rect 5080 245 5126 264
rect 5186 540 5197 586
rect 5243 540 5254 586
rect 5186 426 5254 540
rect 5661 527 5707 549
rect 5865 595 5911 606
rect 5186 425 5806 426
rect 5186 379 5749 425
rect 5795 379 5806 425
rect 4962 172 4973 218
rect 5019 172 5030 218
rect 5186 218 5254 379
rect 5865 368 5911 549
rect 6426 685 6472 724
rect 6009 527 6055 549
rect 6103 549 6213 595
rect 6259 549 6306 595
rect 6103 466 6306 549
rect 6426 527 6472 545
rect 5865 357 6155 368
rect 5865 326 6109 357
rect 5490 280 5501 326
rect 5547 311 6109 326
rect 5547 300 6155 311
rect 5547 280 5910 300
rect 5186 172 5197 218
rect 5243 172 5254 218
rect 5633 210 5679 221
rect 3957 106 4415 152
rect 3722 60 3796 97
rect 4694 71 4705 117
rect 4751 71 4762 117
rect 4694 60 4762 71
rect 5633 60 5679 164
rect 5857 210 5910 280
rect 5903 164 5910 210
rect 5857 151 5910 164
rect 6021 167 6067 178
rect 6021 60 6067 121
rect 6230 167 6306 466
rect 6230 121 6245 167
rect 6291 121 6306 167
rect 6230 110 6306 121
rect 6469 158 6515 178
rect 6469 60 6515 112
rect 0 21 6720 60
rect 0 -31 4075 21
rect 4127 -31 6720 21
rect 0 -60 6720 -31
<< via1 >>
rect 1368 632 1373 678
rect 1373 632 1419 678
rect 1419 632 1420 678
rect 1368 626 1420 632
rect 3958 626 4010 678
rect 1339 106 1391 158
rect 4062 265 4108 306
rect 4108 265 4114 306
rect 4062 254 4114 265
rect 3905 106 3957 158
rect 4075 -31 4127 21
<< metal2 >>
rect 1356 678 4033 683
rect 1356 626 1368 678
rect 1420 627 3958 678
rect 1420 626 1432 627
rect 1356 624 1432 626
rect 3946 626 3958 627
rect 4010 626 4033 678
rect 3946 624 4033 626
rect 4049 310 4131 319
rect 4049 254 4062 310
rect 4118 254 4131 310
rect 4049 243 4131 254
rect 1327 158 1393 160
rect 3893 158 3969 162
rect 1327 106 1339 158
rect 1391 106 3905 158
rect 3957 106 3969 158
rect 1327 102 3960 106
rect 4059 25 4141 33
rect 4059 -31 4075 25
rect 4131 -31 4141 25
rect 4059 -43 4141 -31
<< via2 >>
rect 4062 306 4118 310
rect 4062 254 4114 306
rect 4114 254 4118 306
rect 4075 21 4131 25
rect 4075 -31 4127 21
rect 4127 -31 4131 21
<< metal3 >>
rect 4049 310 4131 321
rect 4049 254 4062 310
rect 4118 254 4131 310
rect 4049 243 4131 254
rect 4068 34 4124 243
rect 4059 25 4141 34
rect 4059 -31 4075 25
rect 4131 -31 4141 25
rect 4059 -43 4141 -31
<< labels >>
flabel metal1 s 0 724 6720 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -60 6720 60 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 3 nsew ground bidirectional
flabel metal1 112 281 240 499 0 FreeSans 600 0 0 0 CLK
port 5 nsew clock input
flabel metal1 3079 466 3282 595 0 FreeSans 600 0 0 0 Q0
port 6 nsew signal output
flabel metal1 1026 242 1107 542 0 FreeSans 600 0 0 0 D0
port 7 nsew signal input
flabel metal1 3206 110 3282 466 0 FreeSans 600 0 0 0 Q0
port 6 nsew signal output
<< end >>
